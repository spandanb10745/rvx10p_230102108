`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: spandan_bharadwaj_230102108
// 
// Create Date: 22.09.2025 07:34:27
// Design Name: 
// Module Name: maindec
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: Main control unit decoder.
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/**
 * @brief Main instruction decoder.
 * @details Uses the 7-bit opcode to generate the primary control signals
 * for the Decode stage.
 *
 * @param op          Input 7-bit instruction opcode.
 * @param ResultSrc   Output signal selecting the data source for write-back.
 * @param MemWrite    Output signal enabling data memory write.
 * @param Branch      Output signal indicating a branch instruction.
 * @param ALUSrc      Output signal selecting the ALU's second operand.
 * @param RegWrite    Output signal enabling register file write.
 * @param Jump        Output signal indicating a jump instruction (JAL).
 * @param ImmSrc      Output signal selecting the immediate format.
 * @param ALUOp       Output 2-bit signal for the ALU decoder.
 */
module maindec(
  input  logic [6:0] op,
  output logic [1:0] ResultSrc,
  output logic       MemWrite,
  output logic       Branch, ALUSrc,
  output logic       RegWrite, Jump,
  output logic [1:0] ImmSrc,
  output logic [1:0] ALUOp
);

  // Internal wire to hold all control signals
  logic [10:0] controls;

  // Assign bits from the 'controls' wire to the respective output ports
  assign {RegWrite, ImmSrc, ALUSrc, MemWrite,
          ResultSrc, Branch, ALUOp, Jump} = controls;

  // Combinational logic to decode the opcode
  always_comb
    case(op)
    //         RegWrite_ImmSrc_ALUSrc_MemWrite_ResultSrc_Branch_ALUOp_Jump
      7'b0000011: controls = 11'b1_00_1_0_01_0_00_0; // lw
      7'b0100011: controls = 11'b0_01_1_1_00_0_00_0; // sw
      7'b0110011: controls = 11'b1_xx_0_0_00_0_10_0; // R-type 
      7'b1100011: controls = 11'b0_10_0_0_00_1_01_0; // beq
      7'b0010011: controls = 11'b1_00_1_0_00_0_10_0; // I-type ALU
      7'b1101111: controls = 11'b1_11_0_0_10_0_00_1; // jal
      7'b0001011: controls = 11'b1_xx_0_0_00_0_11_0; // R-type_newly_added_instructions (RVX10)
      default:    controls = 11'bx_xx_x_x_xx_x_xx_x; // non-implemented instruction
    endcase
endmodule
